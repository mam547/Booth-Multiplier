*
* .CONNECT statements
*
.CONNECT GND 0


* ELDO netlist generated with ICnet by 'gota' on Thu Mar  3 2022 at 19:08:02

*
* Globals.
*
.global GND VDD

*
* Component pathname : $ADK/parts/buf02
*
.subckt BUF02  A Y

        M_I$614 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$615 Y N$411 GND GND n L=0.6u W=3u
        M_I$411 N$411 A VDD VDD p L=0.6u W=2.7u
        M_I$412 N$411 A GND GND n L=0.6u W=1.5u
.ends BUF02

*
* Component pathname : $ADK/parts/inv02
*
.subckt INV02  A Y

        M_I$6 Y A VDD VDD p L=0.6u W=5.4u
        M_I$5 Y A GND GND n L=0.6u W=3u
.ends INV02

*
* Component pathname : $ADK/parts/xor2
*
.subckt XOR2  Y A0 A1

        M_I$421 Y N$4 GND GND n L=0.6u W=1.5u
        M_I$420 Y N$4 VDD VDD p L=0.6u W=2.7u
        M_I$218 N$213 A1 GND GND n L=0.6u W=3u
        M_I$217 N$212 A0 N$213 GND n L=0.6u W=3u
        M_I$9 N$212 A1 VDD VDD p L=0.6u W=3.9u
        M_I$8 N$212 A0 VDD VDD p L=0.6u W=3.9u
        M_I$7 N$3 N$212 GND GND n L=0.6u W=3u
        M_I$6 N$4 A1 N$3 GND n L=0.6u W=3u
        M_I$5 N$4 A0 N$3 GND n L=0.6u W=3u
        M_I$4 N$4 A1 N$1 VDD p L=0.6u W=7.8u
        M_I$3 N$4 N$212 VDD VDD p L=0.6u W=3.9u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=7.8u
.ends XOR2

*
* Component pathname : $ADK/parts/nor02_2x
*
.subckt NOR02_2X  A0 A1 Y

        M_I$5 Y A0 GND GND n L=0.6u W=3u
        M_I$4 Y A1 GND GND n L=0.6u W=3u
        M_I$3 Y A1 N$1 VDD p L=0.6u W=7.8u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=7.8u
.ends NOR02_2X

*
* Component pathname : $ADK/parts/nand02_2x
*
.subckt NAND02_2X  Y A0 A1

        M_I$9 Y A1 VDD VDD p L=0.6u W=6u
        M_I$8 Y A0 VDD VDD p L=0.6u W=6u
        M_I$3 Y A0 N$5 GND n L=0.6u W=6u
        M_I$2 N$5 A1 GND GND n L=0.6u W=6u
.ends NAND02_2X

*
* Component pathname : $ADK/parts/xnor2
*
.subckt XNOR2  Y A0 A1

        M_I$218 N$213 A1 GND GND n L=0.6u W=3u
        M_I$217 N$212 A0 N$213 GND n L=0.6u W=3u
        M_I$9 N$212 A1 VDD VDD p L=0.6u W=3.9u
        M_I$8 N$212 A0 VDD VDD p L=0.6u W=3.9u
        M_I$7 N$3 N$212 GND GND n L=0.6u W=3u
        M_I$6 Y A1 N$3 GND n L=0.6u W=3u
        M_I$5 Y A0 N$3 GND n L=0.6u W=3u
        M_I$4 Y A1 N$1 VDD p L=0.6u W=7.8u
        M_I$3 Y N$212 VDD VDD p L=0.6u W=3.9u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=7.8u
.ends XNOR2

*
* Component pathname : $ADK/parts/nor02ii
*
.subckt NOR02II  A0 A1 Y

        MP1 N$208 A1 VDD VDD p L=0.6u W=2.7u
        MN1 N$208 A1 GND GND n L=0.6u W=1.5u
        MN4 Y A0 GND GND n L=0.6u W=1.5u
        MN2 Y N$208 GND GND n L=0.6u W=1.5u
        MP4 Y N$208 N$4 VDD p L=0.6u W=3.9u
        MP2 N$4 A0 VDD VDD p L=0.6u W=3.9u
.ends NOR02II

*
* Component pathname : $ADK/parts/aoi22
*
.subckt AOI22  B1 A0 A1 B0 Y

        M_I$425 Y B0 N$9 GND n L=0.6u W=3u
        M_I$426 Y B1 N$4 VDD p L=0.6u W=3.9u
        M_I$12 N$8 A1 GND GND n L=0.6u W=3u
        M_I$11 Y A0 N$8 GND n L=0.6u W=3u
        M_I$7 Y B0 N$4 VDD p L=0.6u W=3.9u
        M_I$6 N$4 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$4 A0 VDD VDD p L=0.6u W=3.9u
        M_I$13 N$9 B1 GND GND n L=0.6u W=3u
.ends AOI22

*
* Component pathname : $ADK/parts/mux21
*
.subckt MUX21  S0 A0 A1 Y

        M_I$5 Y S0 N$10 VDD p L=0.6u W=5.4u
        M_I$13 N$6 A1 GND GND n L=0.6u W=3u
        M_I$12 Y S0 N$6 GND n L=0.6u W=3u
        M_I$17 Y N$7 N$5 VDD p L=0.6u W=5.4u
        M_I$16 N$5 A1 VDD VDD p L=0.6u W=5.4u
        M_I$7 N$4 A0 GND GND n L=0.6u W=3u
        M_I$6 Y N$7 N$4 GND n L=0.6u W=3u
        M_I$4 N$10 A0 VDD VDD p L=0.6u W=5.4u
        M_I$3 N$7 S0 GND GND n L=0.6u W=1.5u
        M_I$2 N$7 S0 VDD VDD p L=0.6u W=2.7u
.ends MUX21

*
* Component pathname : $ADK/parts/mux21_ni
*
.subckt MUX21_NI  S0 A0 A1 Y

        M_I$18 Y N$11 GND GND n L=0.6u W=1.5u
        M_I$17 Y N$11 VDD VDD p L=0.6u W=2.7u
        M_I$16 N$11 S0 N$7 VDD p L=0.6u W=5.4u
        M_I$11 N$3 A1 GND GND n L=0.6u W=3u
        M_I$10 N$11 S0 N$3 GND n L=0.6u W=3u
        M_I$9 N$11 N$4 N$2 VDD p L=0.6u W=5.4u
        M_I$8 N$2 A1 VDD VDD p L=0.6u W=5.4u
        M_I$7 N$1 A0 GND GND n L=0.6u W=3u
        M_I$6 N$11 N$4 N$1 GND n L=0.6u W=3u
        M_I$4 N$7 A0 VDD VDD p L=0.6u W=5.4u
        M_I$3 N$4 S0 GND GND n L=0.6u W=1.5u
        M_I$2 N$4 S0 VDD VDD p L=0.6u W=2.7u
.ends MUX21_NI

*
* Component pathname : $ADK/parts/dff
*
.subckt DFF  QB Q CLK D

        M_I$441 N$847 BCLK- N$851 GND n L=0.6u W=4.5u
        M_I$440 N$849 N$847 VDD VDD p L=0.6u W=1.5u
        M_I$439 N$847 BCLK- N$848 VDD p L=0.6u W=1.5u
        M_I$438 N$848 N$849 VDD VDD p L=0.6u W=1.5u
        M_I$437 N$847 BCLK N$845 VDD p L=0.6u W=8.1u
        M_I$436 N$845 D VDD VDD p L=0.6u W=8.1u
        M_I$452 BCLK BCLK- GND GND n L=0.6u W=3u
        M_I$673 Q QB GND GND n L=0.6u W=3u
        M_I$672 Q QB VDD VDD p L=0.6u W=5.4u
        M_I$669 QB N$1074 GND GND n L=0.6u W=3u
        M_I$675 QB N$1074 VDD VDD p L=0.6u W=5.4u
        M_I$668 N$1071 N$1074 GND GND n L=0.6u W=1.5u
        M_I$667 N$1073 N$1071 GND GND n L=0.6u W=1.5u
        M_I$666 N$1074 BCLK- N$1073 GND n L=0.6u W=1.5u
        M_I$665 N$1072 N$847 GND GND n L=0.6u W=4.5u
        M_I$664 N$1074 BCLK N$1072 GND n L=0.6u W=4.5u
        M_I$663 N$1071 N$1074 VDD VDD p L=0.6u W=1.5u
        M_I$662 N$1074 BCLK N$1070 VDD p L=0.6u W=1.5u
        M_I$661 N$1070 N$1071 VDD VDD p L=0.6u W=1.5u
        M_I$660 N$1074 BCLK- N$1069 VDD p L=0.6u W=8.1u
        M_I$659 N$1069 N$847 VDD VDD p L=0.6u W=8.1u
        M_I$449 BCLK- CLK GND GND n L=0.6u W=3u
        M_I$448 BCLK- CLK VDD VDD p L=0.6u W=5.4u
        M_I$453 BCLK BCLK- VDD VDD p L=0.6u W=5.4u
        M_I$445 N$849 N$847 GND GND n L=0.6u W=1.5u
        M_I$444 N$852 N$849 GND GND n L=0.6u W=1.5u
        M_I$443 N$847 BCLK N$852 GND n L=0.6u W=1.5u
        M_I$442 N$851 D GND GND n L=0.6u W=4.5u
.ends DFF

*
* Component pathname : $ADK/parts/oai21
*
.subckt OAI21  A0 A1 B0 Y

        M_I$5 N$7 B0 GND GND n L=0.6u W=3u
        M_I$4 Y A1 N$7 GND n L=0.6u W=3u
        M_I$3 Y A0 N$7 GND n L=0.6u W=3u
        M_I$12 Y B0 VDD VDD p L=0.6u W=3.6u
        M_I$2 Y A1 N$9 VDD p L=0.6u W=7.2u
        M_I$1 N$9 A0 VDD VDD p L=0.6u W=7.2u
.ends OAI21

*
* Component pathname : $ADK/parts/and02
*
.subckt AND02  Y A0 A1

        M_I$674 Y N$5 VDD VDD p L=0.6u W=2.7u
        M_I$675 Y N$5 GND GND n L=0.6u W=1.5u
        M_I$472 N$5 A1 VDD VDD p L=0.6u W=3.6u
        M_I$471 N$5 A0 VDD VDD p L=0.6u W=3.6u
        M_I$4 N$5 A0 N$7 GND n L=0.6u W=3u
        M_I$5 N$7 A1 GND GND n L=0.6u W=3u
.ends AND02

*
* Component pathname : $ADK/parts/or02
*
.subckt OR02  A0 A1 Y

        M_I$212 Y N$5 GND GND n L=0.6u W=1.5u
        M_I$211 Y N$5 VDD VDD p L=0.6u W=2.7u
        M_I$5 N$5 A0 GND GND n L=0.6u W=1.5u
        M_I$4 N$5 A1 GND GND n L=0.6u W=1.5u
        M_I$3 N$5 A1 N$1 VDD p L=0.6u W=3.9u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=3.9u
.ends OR02

*
* Component pathname : $ADK/parts/ao32
*
.subckt AO32  Y A0 A1 A2 B0 B1

        M_I$222 Y N$214 GND GND n L=0.6u W=1.5u
        M_I$221 Y N$214 VDD VDD p L=0.6u W=2.7u
        M_I$12 N$6 B1 GND GND n L=0.6u W=3u
        M_I$11 N$214 B0 N$6 GND n L=0.6u W=3u
        M_I$10 N$5 A2 GND GND n L=0.6u W=4.5u
        M_I$9 N$4 A1 N$5 GND n L=0.6u W=4.5u
        M_I$8 N$214 A0 N$4 GND n L=0.6u W=4.5u
        M_I$6 N$214 B0 N$11 VDD p L=0.6u W=3.9u
        M_I$5 N$214 B1 N$11 VDD p L=0.6u W=3.9u
        M_I$4 N$11 A0 VDD VDD p L=0.6u W=3.9u
        M_I$3 N$11 A1 VDD VDD p L=0.6u W=3.9u
        M_I$2 N$11 A2 VDD VDD p L=0.6u W=3.9u
.ends AO32

*
* Component pathname : $ADK/parts/aoi21
*
.subckt AOI21  A0 A1 B0 Y

        M_I$12 N$8 A1 GND GND n L=0.6u W=3u
        M_I$11 Y A0 N$8 GND n L=0.6u W=3u
        M_I$7 Y B0 N$4 VDD p L=0.6u W=3.9u
        M_I$6 N$4 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$4 A0 VDD VDD p L=0.6u W=3.9u
        M_I$13 Y B0 GND GND n L=0.6u W=1.5u
.ends AOI21

*
* Component pathname : $ADK/parts/nor03
*
.subckt NOR03  A2 A0 A1 Y

        M_I$213 Y A0 GND GND n L=0.6u W=1.8u
        M_I$211 Y A2 N$211 VDD p L=0.6u W=8.1u
        M_I$5 Y A1 GND GND n L=0.6u W=1.8u
        M_I$4 Y A2 GND GND n L=0.6u W=1.8u
        M_I$3 N$211 A1 N$1 VDD p L=0.6u W=8.1u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=8.1u
.ends NOR03

*
* Component pathname : $ADK/parts/nor03_2x
*
.subckt NOR03_2X  A1 A0 A2 Y

        M_I$12 Y A0 GND GND n L=0.6u W=3.3u
        M_I$10 Y A2 N$3 VDD p L=0.6u W=12u
        M_I$5 Y A1 GND GND n L=0.6u W=3.3u
        M_I$4 Y A2 GND GND n L=0.6u W=3.3u
        M_I$3 N$3 A1 N$1 VDD p L=0.6u W=12u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=12u
.ends NOR03_2X

*
* Component pathname : $ADK/parts/aoi221
*
.subckt AOI221  A0 A1 B0 B1 C0 Y

        M_I$13 Y C0 GND GND n L=0.6u W=3u
        M_I$12 N$8 B1 GND GND n L=0.6u W=4.5u
        M_I$11 Y B0 N$8 GND n L=0.6u W=4.5u
        M_I$9 N$6 A1 GND GND n L=0.6u W=4.5u
        M_I$8 Y A0 N$6 GND n L=0.6u W=4.5u
        M_I$7 Y C0 N$4 VDD p L=0.6u W=7.2u
        M_I$6 N$4 B0 N$14 VDD p L=0.6u W=7.2u
        M_I$5 N$4 B1 N$14 VDD p L=0.6u W=7.2u
        M_I$3 N$14 A1 VDD VDD p L=0.6u W=7.2u
        M_I$2 N$14 A0 VDD VDD p L=0.6u W=7.2u
.ends AOI221

*
* Component pathname : $ADK/parts/ao21
*
.subckt AO21  A1 A0 B0 Y

        M_I$14 Y N$3 VDD VDD p L=0.6u W=2.7u
        M_I$13 Y N$3 GND GND n L=0.6u W=1.5u
        M_I$12 N$2 A1 GND GND n L=0.6u W=3u
        M_I$11 N$3 A0 N$2 GND n L=0.6u W=3u
        M_I$7 N$3 B0 N$1 VDD p L=0.6u W=3.9u
        M_I$6 N$1 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$1 A0 VDD VDD p L=0.6u W=3.9u
        M_I$4 N$3 B0 GND GND n L=0.6u W=1.5u
.ends AO21

*
* Component pathname : $ADK/parts/nor04
*
.subckt NOR04  A3 A2 A0 A1 Y

        M_I$415 Y A3 GND GND n L=0.6u W=3u
        M_I$416 Y A3 N$418 VDD p L=0.6u W=10.8u
        M_I$213 Y A0 GND GND n L=0.6u W=3u
        M_I$211 N$418 A2 N$211 VDD p L=0.6u W=10.8u
        M_I$5 Y A1 GND GND n L=0.6u W=3u
        M_I$4 Y A2 GND GND n L=0.6u W=3u
        M_I$3 N$211 A1 N$1 VDD p L=0.6u W=10.8u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=10.8u
.ends NOR04

*
* Component pathname : $ADK/parts/ao22
*
.subckt AO22  A1 A0 B0 Y B1

        M_I$16 Y N$215 VDD VDD p L=0.6u W=2.7u
        M_I$18 Y N$215 GND GND n L=0.6u W=1.5u
        M_I$14 N$215 B0 N$2 GND n L=0.6u W=3u
        M_I$13 N$215 B1 N$6 VDD p L=0.6u W=3.9u
        M_I$12 N$1 A1 GND GND n L=0.6u W=3u
        M_I$11 N$215 A0 N$1 GND n L=0.6u W=3u
        M_I$7 N$215 B0 N$6 VDD p L=0.6u W=3.9u
        M_I$6 N$6 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$6 A0 VDD VDD p L=0.6u W=3.9u
        M_I$4 N$2 B1 GND GND n L=0.6u W=3u
.ends AO22

*
* Component pathname : /home/gota/EECS301/lab3/Multiplier_V/Multiplier_S/Multiplier
*
.subckt MULTIPLIER  MULTIPLICAND[0] MULTIPLICAND[1] MULTIPLICAND[2] MULTIPLICAND[3]
+ MULTIPLIER[0] MULTIPLIER[1] MULTIPLIER[2] MULTIPLIER[3] RESULT[0] RESULT[1]
+ RESULT[2] RESULT[3] RESULT[4] RESULT[5] RESULT[6] RESULT[7] CLK FINISHED
+ START

        X_CL0_IX417 CL0_NX371 CL0_NX418 BUF02
        X_CL0_IX415 CL0_NX313 CL0_NX416 BUF02
        X_CL0_IX409 CL0_NX298 CL0_NX410 INV02
        X_IX548 CL0_NX298 NX549 INV02
        X_CL0_IX161 CL0_NX392 CL0_NX160 INV02
        X_CL0_IX15 CL0_NX362 CL0_NX14 INV02
        X_CL0_IX411 CL0_NX367 CL0_NX412 INV02
        X_CL0_IX299 CL0_NX145 CL0_NX298 INV02
        X_CL0_IX63 CL0_NX321 CL0_NX147 INV02
        X_CL0_IX352 CL0_NX156 M_QREGOUT_0 CL0_M_QNEG XOR2
        X_CL0_IX335 CL0_M_CNT_0 CL0_M_CNT_1 CL0_NX334 NOR02_2X
        X_CL0_IX191 CL0_NX349 CL0_NX367 CL0_NX304 NOR02_2X
        X_CL0_IX393 CL0_NX392 CL0_NX418 CL0_NX156 NAND02_2X
        X_IX169 NX168 NX369 NX166 XNOR2
        X_IX167 NX166 M_ADDSUBA_2 NX164 XNOR2
        X_IX165 NX164 M_ADDSUBCTRL M_ADDSUBB_2 XNOR2
        X_IX225 NX224 M_ADDSUBCTRL M_ADDSUBB_3 XNOR2
        X_IX227 NX226 M_ADDSUBA_3 NX224 XNOR2
        X_IX229 NX228 NX358 NX226 XNOR2
        X_CL0_IX356 CL0_NX416 CL0_NX102 CL0_NX355 NOR02II
        X_CL0_IX101 START CL0_M_NEXTSTATE_2 CL0_NX145 NOR02II
        X_CL0_IX370 CL0_NX319 CL0_NX416 CL0_NX321 CL0_NX418 CL0_NX369 AOI22
        X_CL0_IX83 NX549 CL0_NX345 CL0_NX362 CL0_NX82 MUX21
        X_CL0_IX216 CL0_NX424 CL0_NX319 CL0_NX317 CL0_NX215 MUX21
        X_IX359 NX166 NX164 NX369 NX358 MUX21_NI
        X_CL0_IX236 CL0_NX426 CL0_NX14 NX545 CL0_NX235 MUX21_NI
        X_CL0_IX256 CL0_NX426 CL0_NX82 M_AREGCTRL_0 CL0_NX255 MUX21_NI
        X_CL0_IX226 CL0_NX424 CL0_NX164 FINISHED CL0_NX225 MUX21_NI
        X_CL0_IX196 CL0_NX424 CL0_NX116 CL0_M_NEXTSTATE_0 CL0_NX195 MUX21_NI
        X_CL0_REG_M_QNEG CL0_NX359 CL0_M_QNEG CL0_NX414 CL0_NX205 DFF
        X_CL0_REG_M_NEXTSTATE_1 CL0_NX317 CL0_M_NEXTSTATE_1 CL0_NX414 CL0_NX215 DFF
        X_CL0_REG_M_NEXTSTATE_0 CL0_NX306 CL0_M_NEXTSTATE_0 CL0_NX414 CL0_NX195 DFF
        X_CL0_IX366 NX549 CL0_NX412 CL0_NX349 CL0_NX365 OAI21
        X_CL0_IX363 CL0_NX362 CL0_NX349 CL0_NX367 AND02
        X_CL0_IX185 START CL0_NX317 CL0_NX367 OR02
        X_CL0_IX127 START CL0_NX306 CL0_NX349 OR02
        X_CL0_IX206 CL0_NX205 M_QREGNEG CL0_NX410 CL0_NX416 CL0_M_QNEG CL0_NX355 AO32
        X_CL0_IX286 CL0_NX285 M_QREGOUT_0 CL0_NX359 CL0_NX418 M_ADDSUBCTRL
+ CL0_NX392 AO32
        X_CL0_IX333 CL0_M_CNT_1 CL0_M_CNT_0 CL0_NX334 CL0_NX332 AOI21
        X_CL0_IX184 CL0_NX365 CL0_NX369 CL0_NX424 CL0_NX183 AOI21
        X_CL0_IX264 CL0_NX349 CL0_NX298 CL0_NX424 CL0_NX263 AOI21
        X_CL0_IX154 CL0_NX14 CL0_M_CNT_0 CL0_NX298 CL0_NX153 NOR03
        X_CL0_IX164 CL0_NX14 CL0_NX298 CL0_NX332 CL0_NX163 NOR03
        X_CL0_IX346 CL0_M_NEXTSTATE_0 START CL0_NX317 CL0_NX345 NOR03_2X
        X_CL0_IX320 CL0_NX416 CL0_NX321 CL0_NX410 CL0_NX345 CL0_NX160 CL0_NX319 AOI221
        X_CL0_IX156 CL0_NX14 CL0_M_CNT_0 CL0_NX153 CL0_NX155 AO21
        X_CL0_IX166 CL0_NX14 CL0_M_CNT_1 CL0_NX163 CL0_NX165 AO21
        X_CL0_IX186 CL0_NX424 CL0_M_NEXTSTATE_2 CL0_NX183 CL0_NX185 AO21
        X_CL0_IX117 CL0_NX147 CL0_NX416 CL0_NX362 CL0_NX116 AO21
        X_CL0_IX266 CL0_NX424 M_AREGCTRL_1 CL0_NX263 CL0_NX265 AO21
        X_CL0_IX165 CL0_NX317 CL0_M_NEXTSTATE_0 CL0_NX298 START CL0_NX164 NOR04
        X_CL0_IX372 CL0_NX306 CL0_M_NEXTSTATE_2 START CL0_M_NEXTSTATE_1
+ CL0_NX371 NOR04
        X_CL0_IX314 CL0_NX306 CL0_NX298 START CL0_M_NEXTSTATE_1 CL0_NX313 NOR04
        X_CL0_IX423 CL0_NX304 CL0_NX424 BUF02
        X_CL0_IX425 CL0_NX304 CL0_NX426 BUF02
        X_IX477 M_AREGCTRL_1 NX478 BUF02
        X_IX479 M_MREGCTRL NX480 BUF02
        X_IX481 M_MREGCTRL NX482 BUF02
        X_IX37 M_AREGCTRL_0 NX478 NX36 NOR02_2X
        X_IX31 NX30 NX476 M_AREGCTRL_0 NAND02_2X
        X_IX336 NX36 NX476 AR0_M_REG_1 M_ADDSUBOUT_0 NX335 AOI22
        X_IX350 NX36 NX476 AR0_M_REG_3 M_ADDSUBOUT_2 NX349 AOI22
        X_IX342 NX36 NX476 AR0_M_REG_2 M_ADDSUBOUT_1 NX341 AOI22
        X_IX283 NX30 NX333 NX335 NX282 MUX21
        X_IX250 NX30 NX333 NX335 NX249 MUX21
        X_IX79 NX30 NX339 NX341 NX78 MUX21
        X_IX240 NX30 NX339 NX341 NX239 MUX21
        X_IX140 NX30 NX347 NX349 NX136 MUX21
        X_IX230 NX30 NX347 NX349 NX229 MUX21
        X_IX305 AR0_M_REG_0 NX476 M_ADDSUBOUT_0 NX304 NX36 AO22
        X_IX180 NX480 MR0_M_REG_0 MULTIPLICAND[0] NX179 MUX21_NI
        X_IX53 NX480 MR0_M_REG_0 MULTIPLICAND[0] NX52 MUX21_NI
        X_IX190 NX480 MR0_M_REG_1 MULTIPLICAND[1] NX189 MUX21_NI
        X_IX99 NX480 MR0_M_REG_1 MULTIPLICAND[1] NX98 MUX21_NI
        X_IX200 NX480 MR0_M_REG_2 MULTIPLICAND[2] NX199 MUX21_NI
        X_IX157 NX480 MR0_M_REG_2 MULTIPLICAND[2] NX156 MUX21_NI
        X_IX210 NX480 MR0_M_REG_3 MULTIPLICAND[3] NX209 MUX21_NI
        X_IX217 NX482 MR0_M_REG_3 MULTIPLICAND[3] NX216 MUX21_NI
        X_IX345 M_QREGCTRL_1 MULTIPLIER[0] QR0_M_REG_1 NX344 MUX21_NI
        X_IX355 M_QREGCTRL_1 MULTIPLIER[0] QR0_M_REG_0 NX354 MUX21_NI
        X_IX335 M_QREGCTRL_1 MULTIPLIER[1] QR0_M_REG_2 NX334 MUX21_NI
        X_IX325 M_QREGCTRL_1 MULTIPLIER[2] QR0_M_REG_3 NX324 MUX21_NI
        X_IX315 M_QREGCTRL_1 MULTIPLIER[3] M_QREGCARRY NX314 MUX21_NI
        X_AR0_REG_M_REG_0 NX333 AR0_M_REG_0 CLK NX249 DFF
        X_AR0_REG_M_REG_1 NX339 AR0_M_REG_1 CLK NX239 DFF
        X_AR0_REG_M_REG_2 NX347 AR0_M_REG_2 CLK NX229 DFF
        X_REG_M_RESULT_4 N$DUMMY_ESC1[31] RESULT[4] CLK M_ADDSUBA_0 DFF
        X_QR0_REG_M_O_3 N$DUMMY_ESC1[30] M_QREGOUT_3 CLK NX428 DFF
        X_REG_M_RESULT_3 N$DUMMY_ESC1[29] RESULT[3] CLK M_QREGOUT_3 DFF
        X_QR0_REG_M_O_2 N$DUMMY_ESC1[28] M_QREGOUT_2 CLK NX408 DFF
        X_REG_M_RESULT_2 N$DUMMY_ESC1[27] RESULT[2] CLK M_QREGOUT_2 DFF
        X_QR0_REG_M_O_1 N$DUMMY_ESC1[26] M_QREGOUT_1 CLK NX388 DFF
        X_REG_M_RESULT_1 N$DUMMY_ESC1[25] RESULT[1] CLK M_QREGOUT_1 DFF
        X_REG_M_RESULT_0 N$DUMMY_ESC1[24] RESULT[0] CLK M_QREGOUT_0 DFF
        X_QR0_REG_M_O_0 N$DUMMY_ESC1[23] M_QREGOUT_0 CLK NX368 DFF
        X_AS0_REG_M_O_0 N$DUMMY_ESC1[22] M_ADDSUBOUT_0 CLK NX292 DFF
        X_AS0_REG_M_O_1 N$DUMMY_ESC1[21] M_ADDSUBOUT_1 CLK NX110 DFF
        X_AS0_REG_M_O_2 N$DUMMY_ESC1[20] M_ADDSUBOUT_2 CLK NX168 DFF
        X_MR0_REG_M_REG_3 N$DUMMY_ESC1[19] MR0_M_REG_3 CLK NX209 DFF
        X_MR0_REG_M_O_3 N$DUMMY_ESC1[18] M_ADDSUBB_3 CLK NX216 DFF
        X_AR0_REG_M_O_3 N$DUMMY_ESC1[17] M_ADDSUBA_3 CLK NX196 DFF
        X_AR0_REG_M_O_2 N$DUMMY_ESC1[16] M_ADDSUBA_2 CLK NX136 DFF
        X_MR0_REG_M_REG_1 N$DUMMY_ESC1[15] MR0_M_REG_1 CLK NX189 DFF
        X_MR0_REG_M_O_1 N$DUMMY_ESC1[14] M_ADDSUBB_1 CLK NX98 DFF
        X_AR0_REG_M_O_1 N$DUMMY_ESC1[13] M_ADDSUBA_1 CLK NX78 DFF
        X_MR0_REG_M_REG_0 N$DUMMY_ESC1[12] MR0_M_REG_0 CLK NX179 DFF
        X_MR0_REG_M_O_0 N$DUMMY_ESC1[11] M_ADDSUBB_0 CLK NX52 DFF
        X_AR0_REG_M_O_0 N$DUMMY_ESC1[10] M_ADDSUBA_0 CLK NX282 DFF
        X_MR0_REG_M_REG_2 N$DUMMY_ESC1[9] MR0_M_REG_2 CLK NX199 DFF
        X_MR0_REG_M_O_2 N$DUMMY_ESC1[8] M_ADDSUBB_2 CLK NX156 DFF
        X_AS0_REG_M_O_3 N$DUMMY_ESC1[7] M_ADDSUBOUT_3 CLK NX228 DFF
        X_AR0_REG_M_REG_3 N$DUMMY_ESC1[6] AR0_M_REG_3 CLK NX219 DFF
        X_AR0_REG_M_SHIFTBIT N$DUMMY_ESC1[5] M_QREGCARRY CLK NX304 DFF
        X_QR0_REG_M_REG_3 N$DUMMY_ESC1[4] QR0_M_REG_3 CLK NX259 DFF
        X_QR0_REG_M_REG_2 N$DUMMY_ESC1[3] QR0_M_REG_2 CLK NX269 DFF
        X_QR0_REG_M_REG_1 N$DUMMY_ESC1[2] QR0_M_REG_1 CLK NX279 DFF
        X_QR0_REG_M_REG_0 N$DUMMY_ESC1[1] QR0_M_REG_0 CLK NX289 DFF
        X_QR0_REG_M_SHIFTBIT N$DUMMY_ESC1[0] M_QREGNEG CLK NX299 DFF
        X_IX107 NX106 M_ADDSUBCTRL M_ADDSUBB_1 XNOR2
        X_IX435 M_QREGCTRL_1 NX545 NX434 NOR02II
        X_IX239 M_AREGCTRL_0 M_ADDSUBOUT_3 NX171 NOR02II
        X_IX370 M_ADDSUBA_1 NX70 NX108 NX395 NX369 AOI22
        X_CL0_IX276 CL0_NX426 CL0_NX357 M_MREGCTRL CL0_NX275 MUX21_NI
        X_CL0_IX246 CL0_NX426 CL0_NX102 M_QREGCTRL_1 CL0_NX245 MUX21_NI
        X_IX220 NX476 NX171 AR0_M_REG_3 NX219 MUX21_NI
        X_IX197 NX476 NX171 AR0_M_REG_3 NX196 MUX21_NI
        X_IX260 NX545 NX314 QR0_M_REG_3 NX259 MUX21_NI
        X_IX429 NX547 NX314 QR0_M_REG_3 NX428 MUX21_NI
        X_IX270 NX545 NX324 QR0_M_REG_2 NX269 MUX21_NI
        X_IX409 NX547 NX324 QR0_M_REG_2 NX408 MUX21_NI
        X_IX280 NX545 NX334 QR0_M_REG_1 NX279 MUX21_NI
        X_IX389 NX547 NX334 QR0_M_REG_1 NX388 MUX21_NI
        X_IX290 NX545 NX344 QR0_M_REG_0 NX289 MUX21_NI
        X_IX369 NX545 NX344 QR0_M_REG_0 NX368 MUX21_NI
        X_IX300 NX434 NX354 M_QREGNEG NX299 MUX21_NI
        X_IX71 M_ADDSUBB_0 M_ADDSUBCTRL M_ADDSUBA_0 NX70 MUX21_NI
        X_CL0_REG_M_MSIGNAL N$DUMMY_ESC1[45] M_MREGCTRL CL0_NOT_CLK CL0_NX275 DFF
        X_CL0_REG_M_ADDSUBSIGNAL N$DUMMY_ESC1[44] M_ADDSUBCTRL CL0_NOT_CLK
+ CL0_NX285 DFF
        X_CL0_REG_M_ASIGNAL_1 N$DUMMY_ESC1[43] M_AREGCTRL_1 CL0_NOT_CLK
+ CL0_NX265 DFF
        X_CL0_REG_M_ASIGNAL_0 N$DUMMY_ESC1[42] M_AREGCTRL_0 CL0_NOT_CLK
+ CL0_NX255 DFF
        X_CL0_REG_M_QSIGNAL_1 N$DUMMY_ESC1[41] M_QREGCTRL_1 CL0_NOT_CLK
+ CL0_NX245 DFF
        X_CL0_REG_M_QSIGNAL_0 N$DUMMY_ESC1[40] M_QREGCTRL_0 CL0_NOT_CLK
+ CL0_NX235 DFF
        X_CL0_REG_M_CNT_2 N$DUMMY_ESC1[39] CL0_M_CNT_2 CL0_NX414 CL0_NX175 DFF
        X_CL0_REG_M_CNT_1 N$DUMMY_ESC1[38] CL0_M_CNT_1 CL0_NX414 CL0_NX165 DFF
        X_CL0_REG_M_CNT_0 N$DUMMY_ESC1[37] CL0_M_CNT_0 CL0_NX414 CL0_NX155 DFF
        X_CL0_REG_M_NEXTSTATE_2 N$DUMMY_ESC1[36] CL0_M_NEXTSTATE_2 CL0_NX414
+ CL0_NX185 DFF
        X_CL0_REG_M_FINISHED N$DUMMY_ESC1[35] FINISHED CL0_NOT_CLK CL0_NX225 DFF
        X_REG_M_RESULT_7 N$DUMMY_ESC1[34] RESULT[7] CLK M_ADDSUBA_3 DFF
        X_REG_M_RESULT_6 N$DUMMY_ESC1[33] RESULT[6] CLK M_ADDSUBA_2 DFF
        X_REG_M_RESULT_5 N$DUMMY_ESC1[32] RESULT[5] CLK M_ADDSUBA_1 DFF
        X_CL0_IX341 CL0_M_CNT_2 CL0_NX148 CL0_NX321 CL0_NX340 AOI21
        X_CL0_IX174 CL0_NX340 CL0_NX410 CL0_NX14 CL0_NX173 AOI21
        X_CL0_IX322 CL0_M_CNT_1 CL0_M_CNT_0 CL0_M_CNT_2 CL0_NX321 NOR03_2X
        X_CL0_IX176 CL0_NX14 CL0_M_CNT_2 CL0_NX173 CL0_NX175 AO21
        X_IX475 M_AREGCTRL_1 NX476 BUF02
        X_IX544 M_QREGCTRL_0 NX545 BUF02
        X_IX546 M_QREGCTRL_0 NX547 BUF02
        X_CL0_IX358 CL0_NX102 CL0_NX357 INV02
        X_CL0_IX45 CL0_NX334 CL0_NX148 INV02
        X_IX396 NX106 NX395 INV02
        X_CL0_IX413 CLK CL0_NX414 INV02
        X_CL0_IX311 CLK CL0_NOT_CLK INV02
        X_IX111 NX110 NX70 NX108 XOR2
        X_IX293 NX292 M_ADDSUBA_0 M_ADDSUBB_0 XOR2
        X_CL0_IX103 CL0_NX102 CL0_NX362 CL0_NX298 NAND02_2X
        X_IX109 NX108 M_ADDSUBA_1 NX106 XNOR2
.ends MULTIPLIER

*
* MAIN CELL: Component pathname : /home/gota/EECS301/lab3/TopModel_Multiplier
*
        X_MULTIPLIER1 B0 B1 B2 B3 A0 A1 A2 A3 R0 R1 R2 R3 R4 R5 R6 R7 CLK
+ FINISHED START MULTIPLIER
*
.end
