* Component: /home/gota/EECS301/lab3/TopModel  Viewpoint: ami05a
.INCLUDE /home/gota/EECS301/lab3/TopModel/ami05a/TopModel_ami05a.spi
.INCLUDE /mgc/adk3_1/technology/ic/models/VDD_5.mod
.INCLUDE /mgc/adk3_1/technology/ic/models/ami05.mod
.PROBE TRAN V(CLK) V(START) V(A3) V(A2) V(A1) V(A0) V(B3) V(B2) V(B1) V(B0)
+ V(FINISHED) V(R7) V(R6) V(R5) V(R4) V(R3) V(R2) V(R1) V(R0)

VFORCE__CLK CLK GND pulse (0 5v 2n 1n 1n 25n 50n)

VFORCE__START START GND pulse (0 5v 2n 1n 1n 50n 5000n)

VFORCE__A3 A3 GND dc 0V

VFORCE__A2 A2 GND dc 0V

VFORCE__A1 A1 GND dc 5V

VFORCE__A0 A0 GND dc 5V

VFORCE__B3 B3 GND dc 0V

VFORCE__B2 B2 GND dc 5V

VFORCE__B1 B1 GND dc 5V

VFORCE__B0 B0 GND dc 5V




.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

.TEMP 27 

.TRAN  0 1000N
