*
* .CONNECT statements
*
.CONNECT GND 0


* ELDO netlist generated with ICnet by 'gota' on Thu Mar  3 2022 at 20:00:12

*
* Globals.
*
.global GND VDD

*
* Component pathname : $ADK/parts/nor02ii
*
.subckt NOR02II  A0 A1 Y

        MP1 N$208 A1 VDD VDD p L=0.6u W=2.7u
        MN1 N$208 A1 GND GND n L=0.6u W=1.5u
        MN4 Y A0 GND GND n L=0.6u W=1.5u
        MN2 Y N$208 GND GND n L=0.6u W=1.5u
        MP4 Y N$208 N$4 VDD p L=0.6u W=3.9u
        MP2 N$4 A0 VDD VDD p L=0.6u W=3.9u
.ends NOR02II

*
* Component pathname : $ADK/parts/mux21_ni
*
.subckt MUX21_NI  S0 A0 A1 Y

        M_I$18 Y N$11 GND GND n L=0.6u W=1.5u
        M_I$17 Y N$11 VDD VDD p L=0.6u W=2.7u
        M_I$16 N$11 S0 N$7 VDD p L=0.6u W=5.4u
        M_I$11 N$3 A1 GND GND n L=0.6u W=3u
        M_I$10 N$11 S0 N$3 GND n L=0.6u W=3u
        M_I$9 N$11 N$4 N$2 VDD p L=0.6u W=5.4u
        M_I$8 N$2 A1 VDD VDD p L=0.6u W=5.4u
        M_I$7 N$1 A0 GND GND n L=0.6u W=3u
        M_I$6 N$11 N$4 N$1 GND n L=0.6u W=3u
        M_I$4 N$7 A0 VDD VDD p L=0.6u W=5.4u
        M_I$3 N$4 S0 GND GND n L=0.6u W=1.5u
        M_I$2 N$4 S0 VDD VDD p L=0.6u W=2.7u
.ends MUX21_NI

*
* Component pathname : $ADK/parts/dff
*
.subckt DFF  QB Q CLK D

        M_I$441 N$847 BCLK- N$851 GND n L=0.6u W=4.5u
        M_I$440 N$849 N$847 VDD VDD p L=0.6u W=1.5u
        M_I$439 N$847 BCLK- N$848 VDD p L=0.6u W=1.5u
        M_I$438 N$848 N$849 VDD VDD p L=0.6u W=1.5u
        M_I$437 N$847 BCLK N$845 VDD p L=0.6u W=8.1u
        M_I$436 N$845 D VDD VDD p L=0.6u W=8.1u
        M_I$452 BCLK BCLK- GND GND n L=0.6u W=3u
        M_I$673 Q QB GND GND n L=0.6u W=3u
        M_I$672 Q QB VDD VDD p L=0.6u W=5.4u
        M_I$669 QB N$1074 GND GND n L=0.6u W=3u
        M_I$675 QB N$1074 VDD VDD p L=0.6u W=5.4u
        M_I$668 N$1071 N$1074 GND GND n L=0.6u W=1.5u
        M_I$667 N$1073 N$1071 GND GND n L=0.6u W=1.5u
        M_I$666 N$1074 BCLK- N$1073 GND n L=0.6u W=1.5u
        M_I$665 N$1072 N$847 GND GND n L=0.6u W=4.5u
        M_I$664 N$1074 BCLK N$1072 GND n L=0.6u W=4.5u
        M_I$663 N$1071 N$1074 VDD VDD p L=0.6u W=1.5u
        M_I$662 N$1074 BCLK N$1070 VDD p L=0.6u W=1.5u
        M_I$661 N$1070 N$1071 VDD VDD p L=0.6u W=1.5u
        M_I$660 N$1074 BCLK- N$1069 VDD p L=0.6u W=8.1u
        M_I$659 N$1069 N$847 VDD VDD p L=0.6u W=8.1u
        M_I$449 BCLK- CLK GND GND n L=0.6u W=3u
        M_I$448 BCLK- CLK VDD VDD p L=0.6u W=5.4u
        M_I$453 BCLK BCLK- VDD VDD p L=0.6u W=5.4u
        M_I$445 N$849 N$847 GND GND n L=0.6u W=1.5u
        M_I$444 N$852 N$849 GND GND n L=0.6u W=1.5u
        M_I$443 N$847 BCLK N$852 GND n L=0.6u W=1.5u
        M_I$442 N$851 D GND GND n L=0.6u W=4.5u
.ends DFF

*
* Component pathname : /home/gota/EECS301/lab3/Qreg_V/Qreg_S/Qreg
*
.subckt QREG  IN[0] IN[1] IN[2] IN[3] CTRL[0] CTRL[1] O[0] O[1] O[2] O[3]
+ CLK SHIFTBIT CARRY

        X_IX239 CTRL[1] CTRL[0] NX238 NOR02II
        X_IX125 CTRL[0] NX28 M_REG_3 NX124 MUX21_NI
        X_IX111 CTRL[0] NX38 M_REG_2 NX110 MUX21_NI
        X_IX97 CTRL[0] NX48 M_REG_1 NX96 MUX21_NI
        X_IX83 CTRL[0] NX58 M_REG_0 NX82 MUX21_NI
        X_IX29 CTRL[1] IN[3] CARRY NX28 MUX21_NI
        X_IX170 CTRL[0] NX28 M_REG_3 NX169 MUX21_NI
        X_IX39 CTRL[1] IN[2] M_REG_3 NX38 MUX21_NI
        X_IX180 CTRL[0] NX38 M_REG_2 NX179 MUX21_NI
        X_IX49 CTRL[1] IN[1] M_REG_2 NX48 MUX21_NI
        X_IX190 CTRL[0] NX48 M_REG_1 NX189 MUX21_NI
        X_IX59 CTRL[1] IN[0] M_REG_1 NX58 MUX21_NI
        X_IX200 CTRL[0] NX58 M_REG_0 NX199 MUX21_NI
        X_IX69 CTRL[1] IN[0] M_REG_0 NX68 MUX21_NI
        X_IX210 NX238 NX68 SHIFTBIT NX209 MUX21_NI
        X_REG_M_O_3 N$DUMMY_ESC1[8] O[3] CLK NX124 DFF
        X_REG_M_O_2 N$DUMMY_ESC1[7] O[2] CLK NX110 DFF
        X_REG_M_O_1 N$DUMMY_ESC1[6] O[1] CLK NX96 DFF
        X_REG_M_O_0 N$DUMMY_ESC1[5] O[0] CLK NX82 DFF
        X_REG_M_REG_3 N$DUMMY_ESC1[4] M_REG_3 CLK NX169 DFF
        X_REG_M_REG_2 N$DUMMY_ESC1[3] M_REG_2 CLK NX179 DFF
        X_REG_M_REG_1 N$DUMMY_ESC1[2] M_REG_1 CLK NX189 DFF
        X_REG_M_REG_0 N$DUMMY_ESC1[1] M_REG_0 CLK NX199 DFF
        X_REG_M_SHIFTBIT N$DUMMY_ESC1[0] SHIFTBIT CLK NX209 DFF
.ends QREG

*
* Component pathname : /home/gota/EECS301/lab3/Mreg_V/Mreg_S/Mreg
*
.subckt MREG  IN[0] IN[1] IN[2] IN[3] O[0] O[1] O[2] O[3] CLK CTRL

        X_IX176 CTRL M_REG_3 IN[3] NX175 MUX21_NI
        X_IX73 CTRL M_REG_3 IN[3] NX72 MUX21_NI
        X_IX166 CTRL M_REG_2 IN[2] NX165 MUX21_NI
        X_IX53 CTRL M_REG_2 IN[2] NX52 MUX21_NI
        X_IX156 CTRL M_REG_1 IN[1] NX155 MUX21_NI
        X_IX33 CTRL M_REG_1 IN[1] NX32 MUX21_NI
        X_IX146 CTRL M_REG_0 IN[0] NX145 MUX21_NI
        X_IX13 CTRL M_REG_0 IN[0] NX12 MUX21_NI
        X_REG_M_REG_3 N$DUMMY_ESC1[7] M_REG_3 CLK NX175 DFF
        X_REG_M_O_3 N$DUMMY_ESC1[6] O[3] CLK NX72 DFF
        X_REG_M_REG_2 N$DUMMY_ESC1[5] M_REG_2 CLK NX165 DFF
        X_REG_M_O_2 N$DUMMY_ESC1[4] O[2] CLK NX52 DFF
        X_REG_M_REG_1 N$DUMMY_ESC1[3] M_REG_1 CLK NX155 DFF
        X_REG_M_O_1 N$DUMMY_ESC1[2] O[1] CLK NX32 DFF
        X_REG_M_REG_0 N$DUMMY_ESC1[1] M_REG_0 CLK NX145 DFF
        X_REG_M_O_0 N$DUMMY_ESC1[0] O[0] CLK NX12 DFF
.ends MREG

*
* Component pathname : $ADK/parts/inv02
*
.subckt INV02  A Y

        M_I$6 Y A VDD VDD p L=0.6u W=5.4u
        M_I$5 Y A GND GND n L=0.6u W=3u
.ends INV02

*
* Component pathname : $ADK/parts/ao21
*
.subckt AO21  A1 A0 B0 Y

        M_I$14 Y N$3 VDD VDD p L=0.6u W=2.7u
        M_I$13 Y N$3 GND GND n L=0.6u W=1.5u
        M_I$12 N$2 A1 GND GND n L=0.6u W=3u
        M_I$11 N$3 A0 N$2 GND n L=0.6u W=3u
        M_I$7 N$3 B0 N$1 VDD p L=0.6u W=3.9u
        M_I$6 N$1 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$1 A0 VDD VDD p L=0.6u W=3.9u
        M_I$4 N$3 B0 GND GND n L=0.6u W=1.5u
.ends AO21

*
* Component pathname : $ADK/parts/nor04
*
.subckt NOR04  A3 A2 A0 A1 Y

        M_I$415 Y A3 GND GND n L=0.6u W=3u
        M_I$416 Y A3 N$418 VDD p L=0.6u W=10.8u
        M_I$213 Y A0 GND GND n L=0.6u W=3u
        M_I$211 N$418 A2 N$211 VDD p L=0.6u W=10.8u
        M_I$5 Y A1 GND GND n L=0.6u W=3u
        M_I$4 Y A2 GND GND n L=0.6u W=3u
        M_I$3 N$211 A1 N$1 VDD p L=0.6u W=10.8u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=10.8u
.ends NOR04

*
* Component pathname : $ADK/parts/mux21
*
.subckt MUX21  S0 A0 A1 Y

        M_I$5 Y S0 N$10 VDD p L=0.6u W=5.4u
        M_I$13 N$6 A1 GND GND n L=0.6u W=3u
        M_I$12 Y S0 N$6 GND n L=0.6u W=3u
        M_I$17 Y N$7 N$5 VDD p L=0.6u W=5.4u
        M_I$16 N$5 A1 VDD VDD p L=0.6u W=5.4u
        M_I$7 N$4 A0 GND GND n L=0.6u W=3u
        M_I$6 Y N$7 N$4 GND n L=0.6u W=3u
        M_I$4 N$10 A0 VDD VDD p L=0.6u W=5.4u
        M_I$3 N$7 S0 GND GND n L=0.6u W=1.5u
        M_I$2 N$7 S0 VDD VDD p L=0.6u W=2.7u
.ends MUX21

*
* Component pathname : $ADK/parts/buf02
*
.subckt BUF02  A Y

        M_I$614 Y N$411 VDD VDD p L=0.6u W=5.4u
        M_I$615 Y N$411 GND GND n L=0.6u W=3u
        M_I$411 N$411 A VDD VDD p L=0.6u W=2.7u
        M_I$412 N$411 A GND GND n L=0.6u W=1.5u
.ends BUF02

*
* Component pathname : $ADK/parts/nand02_2x
*
.subckt NAND02_2X  Y A0 A1

        M_I$9 Y A1 VDD VDD p L=0.6u W=6u
        M_I$8 Y A0 VDD VDD p L=0.6u W=6u
        M_I$3 Y A0 N$5 GND n L=0.6u W=6u
        M_I$2 N$5 A1 GND GND n L=0.6u W=6u
.ends NAND02_2X

*
* Component pathname : $ADK/parts/aoi22
*
.subckt AOI22  B1 A0 A1 B0 Y

        M_I$425 Y B0 N$9 GND n L=0.6u W=3u
        M_I$426 Y B1 N$4 VDD p L=0.6u W=3.9u
        M_I$12 N$8 A1 GND GND n L=0.6u W=3u
        M_I$11 Y A0 N$8 GND n L=0.6u W=3u
        M_I$7 Y B0 N$4 VDD p L=0.6u W=3.9u
        M_I$6 N$4 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$4 A0 VDD VDD p L=0.6u W=3.9u
        M_I$13 N$9 B1 GND GND n L=0.6u W=3u
.ends AOI22

*
* Component pathname : $ADK/parts/ao32
*
.subckt AO32  Y A0 A1 A2 B0 B1

        M_I$222 Y N$214 GND GND n L=0.6u W=1.5u
        M_I$221 Y N$214 VDD VDD p L=0.6u W=2.7u
        M_I$12 N$6 B1 GND GND n L=0.6u W=3u
        M_I$11 N$214 B0 N$6 GND n L=0.6u W=3u
        M_I$10 N$5 A2 GND GND n L=0.6u W=4.5u
        M_I$9 N$4 A1 N$5 GND n L=0.6u W=4.5u
        M_I$8 N$214 A0 N$4 GND n L=0.6u W=4.5u
        M_I$6 N$214 B0 N$11 VDD p L=0.6u W=3.9u
        M_I$5 N$214 B1 N$11 VDD p L=0.6u W=3.9u
        M_I$4 N$11 A0 VDD VDD p L=0.6u W=3.9u
        M_I$3 N$11 A1 VDD VDD p L=0.6u W=3.9u
        M_I$2 N$11 A2 VDD VDD p L=0.6u W=3.9u
.ends AO32

*
* Component pathname : $ADK/parts/nor02_2x
*
.subckt NOR02_2X  A0 A1 Y

        M_I$5 Y A0 GND GND n L=0.6u W=3u
        M_I$4 Y A1 GND GND n L=0.6u W=3u
        M_I$3 Y A1 N$1 VDD p L=0.6u W=7.8u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=7.8u
.ends NOR02_2X

*
* Component pathname : $ADK/parts/aoi21
*
.subckt AOI21  A0 A1 B0 Y

        M_I$12 N$8 A1 GND GND n L=0.6u W=3u
        M_I$11 Y A0 N$8 GND n L=0.6u W=3u
        M_I$7 Y B0 N$4 VDD p L=0.6u W=3.9u
        M_I$6 N$4 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$4 A0 VDD VDD p L=0.6u W=3.9u
        M_I$13 Y B0 GND GND n L=0.6u W=1.5u
.ends AOI21

*
* Component pathname : $ADK/parts/nor03
*
.subckt NOR03  A2 A0 A1 Y

        M_I$213 Y A0 GND GND n L=0.6u W=1.8u
        M_I$211 Y A2 N$211 VDD p L=0.6u W=8.1u
        M_I$5 Y A1 GND GND n L=0.6u W=1.8u
        M_I$4 Y A2 GND GND n L=0.6u W=1.8u
        M_I$3 N$211 A1 N$1 VDD p L=0.6u W=8.1u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=8.1u
.ends NOR03

*
* Component pathname : $ADK/parts/nor03_2x
*
.subckt NOR03_2X  A1 A0 A2 Y

        M_I$12 Y A0 GND GND n L=0.6u W=3.3u
        M_I$10 Y A2 N$3 VDD p L=0.6u W=12u
        M_I$5 Y A1 GND GND n L=0.6u W=3.3u
        M_I$4 Y A2 GND GND n L=0.6u W=3.3u
        M_I$3 N$3 A1 N$1 VDD p L=0.6u W=12u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=12u
.ends NOR03_2X

*
* Component pathname : $ADK/parts/aoi221
*
.subckt AOI221  A0 A1 B0 B1 C0 Y

        M_I$13 Y C0 GND GND n L=0.6u W=3u
        M_I$12 N$8 B1 GND GND n L=0.6u W=4.5u
        M_I$11 Y B0 N$8 GND n L=0.6u W=4.5u
        M_I$9 N$6 A1 GND GND n L=0.6u W=4.5u
        M_I$8 Y A0 N$6 GND n L=0.6u W=4.5u
        M_I$7 Y C0 N$4 VDD p L=0.6u W=7.2u
        M_I$6 N$4 B0 N$14 VDD p L=0.6u W=7.2u
        M_I$5 N$4 B1 N$14 VDD p L=0.6u W=7.2u
        M_I$3 N$14 A1 VDD VDD p L=0.6u W=7.2u
        M_I$2 N$14 A0 VDD VDD p L=0.6u W=7.2u
.ends AOI221

*
* Component pathname : $ADK/parts/oai21
*
.subckt OAI21  A0 A1 B0 Y

        M_I$5 N$7 B0 GND GND n L=0.6u W=3u
        M_I$4 Y A1 N$7 GND n L=0.6u W=3u
        M_I$3 Y A0 N$7 GND n L=0.6u W=3u
        M_I$12 Y B0 VDD VDD p L=0.6u W=3.6u
        M_I$2 Y A1 N$9 VDD p L=0.6u W=7.2u
        M_I$1 N$9 A0 VDD VDD p L=0.6u W=7.2u
.ends OAI21

*
* Component pathname : $ADK/parts/and02
*
.subckt AND02  Y A0 A1

        M_I$674 Y N$5 VDD VDD p L=0.6u W=2.7u
        M_I$675 Y N$5 GND GND n L=0.6u W=1.5u
        M_I$472 N$5 A1 VDD VDD p L=0.6u W=3.6u
        M_I$471 N$5 A0 VDD VDD p L=0.6u W=3.6u
        M_I$4 N$5 A0 N$7 GND n L=0.6u W=3u
        M_I$5 N$7 A1 GND GND n L=0.6u W=3u
.ends AND02

*
* Component pathname : $ADK/parts/xnor2
*
.subckt XNOR2  Y A0 A1

        M_I$218 N$213 A1 GND GND n L=0.6u W=3u
        M_I$217 N$212 A0 N$213 GND n L=0.6u W=3u
        M_I$9 N$212 A1 VDD VDD p L=0.6u W=3.9u
        M_I$8 N$212 A0 VDD VDD p L=0.6u W=3.9u
        M_I$7 N$3 N$212 GND GND n L=0.6u W=3u
        M_I$6 Y A1 N$3 GND n L=0.6u W=3u
        M_I$5 Y A0 N$3 GND n L=0.6u W=3u
        M_I$4 Y A1 N$1 VDD p L=0.6u W=7.8u
        M_I$3 Y N$212 VDD VDD p L=0.6u W=3.9u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=7.8u
.ends XNOR2

*
* Component pathname : $ADK/parts/or02
*
.subckt OR02  A0 A1 Y

        M_I$212 Y N$5 GND GND n L=0.6u W=1.5u
        M_I$211 Y N$5 VDD VDD p L=0.6u W=2.7u
        M_I$5 N$5 A0 GND GND n L=0.6u W=1.5u
        M_I$4 N$5 A1 GND GND n L=0.6u W=1.5u
        M_I$3 N$5 A1 N$1 VDD p L=0.6u W=3.9u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=3.9u
.ends OR02

*
* Component pathname : /home/gota/EECS301/lab3/Control_V/Control_S/ControlLogic
*
.subckt CONTROLLOGIC  QREG[0] QREG[1] QREG[2] QREG[3] ASIGNAL[0] ASIGNAL[1]
+ QSIGNAL[0] QSIGNAL[1] CLK FINISHED ADDSUBSIGNAL MSIGNAL START QNEG

        X_IX706 NX662 NX707 INV02
        X_IX704 NX593 NX705 INV02
        X_IX594 NX440 NX593 INV02
        X_IX15 NX657 NX14 INV02
        X_IX63 NX616 NX442 INV02
        X_IX45 NX629 NX443 INV02
        X_IX653 NX102 NX652 INV02
        X_IX161 NX687 NX160 INV02
        X_IX606 CLK NOT_CLK INV02
        X_IX561 NX719 ASIGNAL[1] NX558 NX560 AO21
        X_IX471 NX14 M_CNT_2 NX468 NX470 AO21
        X_IX461 NX14 M_CNT_1 NX458 NX460 AO21
        X_IX451 NX14 M_CNT_0 NX448 NX450 AO21
        X_IX117 NX442 NX711 NX657 NX116 AO21
        X_IX481 NX719 M_NEXTSTATE_2 NX478 NX480 AO21
        X_IX667 NX601 M_NEXTSTATE_2 START M_NEXTSTATE_1 NX666 NOR04
        X_IX609 NX601 NX593 START M_NEXTSTATE_1 NX608 NOR04
        X_IX165 NX612 M_NEXTSTATE_0 NX593 START NX164 NOR04
        X_REG_M_MSIGNAL N$DUMMY_ESC1[10] MSIGNAL NOT_CLK NX570 DFF
        X_REG_M_ADDSUBSIGNAL N$DUMMY_ESC1[9] ADDSUBSIGNAL NOT_CLK NX580 DFF
        X_REG_M_ASIGNAL_1 N$DUMMY_ESC1[8] ASIGNAL[1] NOT_CLK NX560 DFF
        X_REG_M_ASIGNAL_0 N$DUMMY_ESC1[7] ASIGNAL[0] NOT_CLK NX550 DFF
        X_REG_M_QSIGNAL_1 N$DUMMY_ESC1[6] QSIGNAL[1] NOT_CLK NX540 DFF
        X_REG_M_QSIGNAL_0 N$DUMMY_ESC1[5] QSIGNAL[0] NOT_CLK NX530 DFF
        X_REG_M_QNEG NX654 M_QNEG NX709 NX500 DFF
        X_REG_M_CNT_2 N$DUMMY_ESC1[4] M_CNT_2 NX709 NX470 DFF
        X_REG_M_CNT_1 N$DUMMY_ESC1[3] M_CNT_1 NX709 NX460 DFF
        X_REG_M_CNT_0 N$DUMMY_ESC1[2] M_CNT_0 NX709 NX450 DFF
        X_REG_M_NEXTSTATE_1 NX612 M_NEXTSTATE_1 NX709 NX510 DFF
        X_REG_M_NEXTSTATE_0 NX601 M_NEXTSTATE_0 NX709 NX490 DFF
        X_REG_M_NEXTSTATE_2 N$DUMMY_ESC1[1] M_NEXTSTATE_2 NX709 NX480 DFF
        X_REG_M_FINISHED N$DUMMY_ESC1[0] FINISHED NOT_CLK NX520 DFF
        X_IX83 NX593 NX657 NX640 NX82 MUX21
        X_IX511 NX719 NX614 NX612 NX510 MUX21
        X_IX571 NX721 NX652 MSIGNAL NX570 MUX21_NI
        X_IX551 NX721 NX82 ASIGNAL[0] NX550 MUX21_NI
        X_IX541 NX721 NX102 QSIGNAL[1] NX540 MUX21_NI
        X_IX531 NX721 NX14 QSIGNAL[0] NX530 MUX21_NI
        X_IX491 NX719 NX116 M_NEXTSTATE_0 NX490 MUX21_NI
        X_IX521 NX719 NX164 FINISHED NX520 MUX21_NI
        X_IX720 NX599 NX721 BUF02
        X_IX718 NX599 NX719 BUF02
        X_IX712 NX666 NX713 BUF02
        X_IX710 NX608 NX711 BUF02
        X_IX688 NX687 NX713 NX156 NAND02_2X
        X_IX103 NX102 NX657 NX593 NAND02_2X
        X_IX665 NX614 NX711 NX616 NX713 NX664 AOI22
        X_IX581 NX580 QREG[0] NX654 NX713 ADDSUBSIGNAL NX687 AO32
        X_IX501 NX500 QNEG NX705 NX711 M_QNEG NX650 AO32
        X_IX651 NX711 NX102 NX650 NOR02II
        X_IX101 START M_NEXTSTATE_2 NX440 NOR02II
        X_IX191 NX644 NX662 NX599 NOR02_2X
        X_IX630 M_CNT_0 M_CNT_1 NX629 NOR02_2X
        X_IX559 NX644 NX593 NX719 NX558 AOI21
        X_IX479 NX660 NX664 NX719 NX478 AOI21
        X_IX636 M_CNT_2 NX443 NX616 NX635 AOI21
        X_IX469 NX635 NX705 NX14 NX468 AOI21
        X_IX628 M_CNT_1 M_CNT_0 NX629 NX627 AOI21
        X_IX459 NX14 NX593 NX627 NX458 NOR03
        X_IX449 NX14 M_CNT_0 NX593 NX448 NOR03
        X_IX641 M_NEXTSTATE_0 START NX612 NX640 NOR03_2X
        X_IX617 M_CNT_1 M_CNT_0 M_CNT_2 NX616 NOR03_2X
        X_IX615 NX711 NX616 NX705 NX640 NX160 NX614 AOI221
        X_IX708 CLK NX709 INV02
        X_IX661 NX440 NX707 NX644 NX660 OAI21
        X_IX658 NX657 NX644 NX662 AND02
        X_IX647 NX156 QREG[0] NX654 XNOR2
        X_IX185 START NX612 NX662 OR02
        X_IX127 START NX601 NX644 OR02
.ends CONTROLLOGIC

*
* Component pathname : $ADK/parts/ao22
*
.subckt AO22  A1 A0 B0 Y B1

        M_I$16 Y N$215 VDD VDD p L=0.6u W=2.7u
        M_I$18 Y N$215 GND GND n L=0.6u W=1.5u
        M_I$14 N$215 B0 N$2 GND n L=0.6u W=3u
        M_I$13 N$215 B1 N$6 VDD p L=0.6u W=3.9u
        M_I$12 N$1 A1 GND GND n L=0.6u W=3u
        M_I$11 N$215 A0 N$1 GND n L=0.6u W=3u
        M_I$7 N$215 B0 N$6 VDD p L=0.6u W=3.9u
        M_I$6 N$6 A1 VDD VDD p L=0.6u W=3.9u
        M_I$5 N$6 A0 VDD VDD p L=0.6u W=3.9u
        M_I$4 N$2 B1 GND GND n L=0.6u W=3u
.ends AO22

*
* Component pathname : /home/gota/EECS301/lab3/Areg_V/Areg_S/Areg
*
.subckt AREG  IN[0] IN[1] IN[2] IN[3] CTRL[0] CTRL[1] O[0] O[1] O[2] O[3]
+ CLK SHIFTBIT

        X_IX13 NX12 CTRL[1] CTRL[0] NAND02_2X
        X_IX5 CTRL[0] CTRL[1] NX4 NOR02_2X
        X_IX25 CTRL[0] IN[3] NX24 NOR02II
        X_IX121 CTRL[1] NX24 M_REG_3 NX120 MUX21_NI
        X_IX140 CTRL[1] NX24 M_REG_3 NX139 MUX21_NI
        X_IX198 NX4 CTRL[1] M_REG_3 IN[2] NX197 AOI22
        X_IX192 NX4 CTRL[1] M_REG_2 IN[1] NX191 AOI22
        X_IX186 NX4 CTRL[1] M_REG_1 IN[0] NX185 AOI22
        X_IX107 NX12 NX195 NX197 NX106 MUX21
        X_IX93 NX12 NX189 NX191 NX92 MUX21
        X_IX79 NX12 NX183 NX185 NX78 MUX21
        X_IX150 NX12 NX195 NX197 NX149 MUX21
        X_IX160 NX12 NX189 NX191 NX159 MUX21
        X_IX170 NX12 NX183 NX185 NX169 MUX21
        X_IX65 M_REG_0 CTRL[1] IN[0] NX64 NX4 AO22
        X_REG_M_O_3 N$DUMMY_ESC1[5] O[3] CLK NX120 DFF
        X_REG_M_O_2 N$DUMMY_ESC1[4] O[2] CLK NX106 DFF
        X_REG_M_O_1 N$DUMMY_ESC1[3] O[1] CLK NX92 DFF
        X_REG_M_O_0 N$DUMMY_ESC1[2] O[0] CLK NX78 DFF
        X_REG_M_REG_3 N$DUMMY_ESC1[1] M_REG_3 CLK NX139 DFF
        X_REG_M_REG_2 NX195 M_REG_2 CLK NX149 DFF
        X_REG_M_REG_1 NX189 M_REG_1 CLK NX159 DFF
        X_REG_M_REG_0 NX183 M_REG_0 CLK NX169 DFF
        X_REG_M_SHIFTBIT N$DUMMY_ESC1[0] SHIFTBIT CLK NX64 DFF
.ends AREG

*
* Component pathname : $ADK/parts/xor2
*
.subckt XOR2  Y A0 A1

        M_I$421 Y N$4 GND GND n L=0.6u W=1.5u
        M_I$420 Y N$4 VDD VDD p L=0.6u W=2.7u
        M_I$218 N$213 A1 GND GND n L=0.6u W=3u
        M_I$217 N$212 A0 N$213 GND n L=0.6u W=3u
        M_I$9 N$212 A1 VDD VDD p L=0.6u W=3.9u
        M_I$8 N$212 A0 VDD VDD p L=0.6u W=3.9u
        M_I$7 N$3 N$212 GND GND n L=0.6u W=3u
        M_I$6 N$4 A1 N$3 GND n L=0.6u W=3u
        M_I$5 N$4 A0 N$3 GND n L=0.6u W=3u
        M_I$4 N$4 A1 N$1 VDD p L=0.6u W=7.8u
        M_I$3 N$4 N$212 VDD VDD p L=0.6u W=3.9u
        M_I$2 N$1 A0 VDD VDD p L=0.6u W=7.8u
.ends XOR2

*
* Component pathname : /home/gota/EECS301/lab3/AddSub_V/AddSub_S/AddSub
*
.subckt ADDSUB  A[0] A[1] A[2] A[3] B[0] B[1] B[2] B[3] O[0] O[1] O[2] O[3]
+ CLK CTRL

        X_IX159 NX22 NX158 INV02
        X_IX157 NX24 NX158 A[1] NX20 NX156 AOI22
        X_IX67 NX66 B[3] CTRL XNOR2
        X_IX69 NX68 A[3] NX66 XNOR2
        X_IX71 NX70 NX167 NX68 XNOR2
        X_IX45 NX44 B[2] CTRL XNOR2
        X_IX47 NX46 A[2] NX44 XNOR2
        X_IX49 NX48 NX156 NX46 XNOR2
        X_IX23 NX22 B[1] CTRL XNOR2
        X_IX25 NX24 A[1] NX22 XNOR2
        X_IX168 NX46 NX44 NX156 NX167 MUX21_NI
        X_IX21 B[0] CTRL A[0] NX20 MUX21_NI
        X_IX27 NX26 NX20 NX24 XOR2
        X_IX5 NX4 A[0] B[0] XOR2
        X_REG_M_O_3 N$DUMMY_ESC1[3] O[3] CLK NX70 DFF
        X_REG_M_O_2 N$DUMMY_ESC1[2] O[2] CLK NX48 DFF
        X_REG_M_O_1 N$DUMMY_ESC1[1] O[1] CLK NX26 DFF
        X_REG_M_O_0 N$DUMMY_ESC1[0] O[0] CLK NX4 DFF
.ends ADDSUB

*
* MAIN CELL: Component pathname : /home/gota/EECS301/lab3/TopModel
*
        X_QREG1 B0 B1 B2 B3 N$35[0] N$35[1] R0 R1 R2 R3 CLK N$33 N$28 QREG
        X_MREG1 A0 A1 A2 A3 N$8[0] N$8[1] N$8[2] N$8[3] CLK N$22 MREG
        X_CONTROLLOGIC1 R0 R1 R2 R3 N$29[0] N$29[1] N$35[0] N$35[1] CLK
+ FINISHED N$48 N$22 START N$33 CONTROLLOGIC
        X_AREG1 N$18[0] N$18[1] N$18[2] N$18[3] N$29[0] N$29[1] R4 R5 R6
+ R7 CLK N$28 AREG
        X_ADDSUB1 R4 R5 R6 R7 N$8[0] N$8[1] N$8[2] N$8[3] N$18[0] N$18[1]
+ N$18[2] N$18[3] CLK N$48 ADDSUB
*
.end
